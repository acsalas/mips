module bcd2seven( bcd, segs);

//input rst;
input [3:0] bcd;
output [6:0] segs;

assign segs =  (bcd == 4'b0000)?7'b1000000:(bcd == 4'b0001)?7'b1111001:(bcd == 4'b0010)?7'b0100100:(bcd == 4'b0011)?7'b0110000:
					(bcd == 4'b0100)?7'b0011001:(bcd == 4'b0101)?7'b0010010:(bcd == 4'b0110)?7'b0000010:(bcd == 4'b0111)?7'b1111000:
					(bcd == 4'b1000)?7'b0000000:(bcd == 4'b1001)?7'b0011000:(bcd == 4'b1010)?7'b0001000:(bcd == 4'b1011)?7'b0000011:
					(bcd == 4'b1100)?7'b1000110:(bcd == 4'b1101)?7'b0100001:(bcd == 4'b1110)?7'b0000110:7'b0001110;
				
				
endmodule
